/escnfs/courses/fa24-cse-30342.01/dropbox/mjohns79/VLSI/lab5solo/muddlib.lef